module tb_uart_tx;

reg i_Clock;
reg i_TX_DV;
reg [7:0] i_TX_Byte;
wire o_TX_Active;
wire o_uart_tx;
wire o_TX_Done;

initial begin
    $from_myhdl(
        i_Clock,
        i_TX_DV,
        i_TX_Byte
    );
    $to_myhdl(
        o_TX_Active,
        o_uart_tx,
        o_TX_Done
    );
end

uart_tx dut(
    i_Clock,
    i_TX_DV,
    i_TX_Byte,
    o_TX_Active,
    o_uart_tx,
    o_TX_Done
);

endmodule
